
module soc_design (
	clock_clk,
	fpga_reset_n);	

	input		clock_clk;
	input		fpga_reset_n;
endmodule
