// hps_design.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module hps_design (
		input  wire        clk_clk,             //         clk.clk
		output wire [14:0] hps_ddr_mem_a,       //     hps_ddr.mem_a
		output wire [2:0]  hps_ddr_mem_ba,      //            .mem_ba
		output wire        hps_ddr_mem_ck,      //            .mem_ck
		output wire        hps_ddr_mem_ck_n,    //            .mem_ck_n
		output wire        hps_ddr_mem_cke,     //            .mem_cke
		output wire        hps_ddr_mem_cs_n,    //            .mem_cs_n
		output wire        hps_ddr_mem_ras_n,   //            .mem_ras_n
		output wire        hps_ddr_mem_cas_n,   //            .mem_cas_n
		output wire        hps_ddr_mem_we_n,    //            .mem_we_n
		output wire        hps_ddr_mem_reset_n, //            .mem_reset_n
		inout  wire [31:0] hps_ddr_mem_dq,      //            .mem_dq
		inout  wire [3:0]  hps_ddr_mem_dqs,     //            .mem_dqs
		inout  wire [3:0]  hps_ddr_mem_dqs_n,   //            .mem_dqs_n
		output wire        hps_ddr_mem_odt,     //            .mem_odt
		output wire [3:0]  hps_ddr_mem_dm,      //            .mem_dm
		input  wire        hps_ddr_oct_rzqin,   //            .oct_rzqin
		output wire        ledr_export,         //        ledr.export
		output wire        pll_0_sdram_clk      // pll_0_sdram.clk
	);

	wire         pll_0_outclk0_clk;                     // pll_0:outclk_0 -> [SMP_HPS:h2f_lw_axi_clk, mm_interconnect_0:pll_0_outclk0_clk, pio_0:clk, rst_controller:clk, rst_controller_001:clk]
	wire         smp_hps_h2f_reset_reset;               // SMP_HPS:h2f_rst_n -> [pll_0:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire   [1:0] smp_hps_h2f_lw_axi_master_awburst;     // SMP_HPS:h2f_lw_AWBURST -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awburst
	wire   [3:0] smp_hps_h2f_lw_axi_master_arlen;       // SMP_HPS:h2f_lw_ARLEN -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_arlen
	wire   [3:0] smp_hps_h2f_lw_axi_master_wstrb;       // SMP_HPS:h2f_lw_WSTRB -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_wstrb
	wire         smp_hps_h2f_lw_axi_master_wready;      // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_wready -> SMP_HPS:h2f_lw_WREADY
	wire  [11:0] smp_hps_h2f_lw_axi_master_rid;         // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_rid -> SMP_HPS:h2f_lw_RID
	wire         smp_hps_h2f_lw_axi_master_rready;      // SMP_HPS:h2f_lw_RREADY -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_rready
	wire   [3:0] smp_hps_h2f_lw_axi_master_awlen;       // SMP_HPS:h2f_lw_AWLEN -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awlen
	wire  [11:0] smp_hps_h2f_lw_axi_master_wid;         // SMP_HPS:h2f_lw_WID -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_wid
	wire   [3:0] smp_hps_h2f_lw_axi_master_arcache;     // SMP_HPS:h2f_lw_ARCACHE -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_arcache
	wire         smp_hps_h2f_lw_axi_master_wvalid;      // SMP_HPS:h2f_lw_WVALID -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_wvalid
	wire  [20:0] smp_hps_h2f_lw_axi_master_araddr;      // SMP_HPS:h2f_lw_ARADDR -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_araddr
	wire   [2:0] smp_hps_h2f_lw_axi_master_arprot;      // SMP_HPS:h2f_lw_ARPROT -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_arprot
	wire   [2:0] smp_hps_h2f_lw_axi_master_awprot;      // SMP_HPS:h2f_lw_AWPROT -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awprot
	wire  [31:0] smp_hps_h2f_lw_axi_master_wdata;       // SMP_HPS:h2f_lw_WDATA -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_wdata
	wire         smp_hps_h2f_lw_axi_master_arvalid;     // SMP_HPS:h2f_lw_ARVALID -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_arvalid
	wire   [3:0] smp_hps_h2f_lw_axi_master_awcache;     // SMP_HPS:h2f_lw_AWCACHE -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awcache
	wire  [11:0] smp_hps_h2f_lw_axi_master_arid;        // SMP_HPS:h2f_lw_ARID -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_arid
	wire   [1:0] smp_hps_h2f_lw_axi_master_arlock;      // SMP_HPS:h2f_lw_ARLOCK -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_arlock
	wire   [1:0] smp_hps_h2f_lw_axi_master_awlock;      // SMP_HPS:h2f_lw_AWLOCK -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awlock
	wire  [20:0] smp_hps_h2f_lw_axi_master_awaddr;      // SMP_HPS:h2f_lw_AWADDR -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awaddr
	wire   [1:0] smp_hps_h2f_lw_axi_master_bresp;       // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_bresp -> SMP_HPS:h2f_lw_BRESP
	wire         smp_hps_h2f_lw_axi_master_arready;     // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_arready -> SMP_HPS:h2f_lw_ARREADY
	wire  [31:0] smp_hps_h2f_lw_axi_master_rdata;       // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_rdata -> SMP_HPS:h2f_lw_RDATA
	wire         smp_hps_h2f_lw_axi_master_awready;     // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awready -> SMP_HPS:h2f_lw_AWREADY
	wire   [1:0] smp_hps_h2f_lw_axi_master_arburst;     // SMP_HPS:h2f_lw_ARBURST -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_arburst
	wire   [2:0] smp_hps_h2f_lw_axi_master_arsize;      // SMP_HPS:h2f_lw_ARSIZE -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_arsize
	wire         smp_hps_h2f_lw_axi_master_bready;      // SMP_HPS:h2f_lw_BREADY -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_bready
	wire         smp_hps_h2f_lw_axi_master_rlast;       // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_rlast -> SMP_HPS:h2f_lw_RLAST
	wire         smp_hps_h2f_lw_axi_master_wlast;       // SMP_HPS:h2f_lw_WLAST -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_wlast
	wire   [1:0] smp_hps_h2f_lw_axi_master_rresp;       // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_rresp -> SMP_HPS:h2f_lw_RRESP
	wire  [11:0] smp_hps_h2f_lw_axi_master_awid;        // SMP_HPS:h2f_lw_AWID -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awid
	wire  [11:0] smp_hps_h2f_lw_axi_master_bid;         // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_bid -> SMP_HPS:h2f_lw_BID
	wire         smp_hps_h2f_lw_axi_master_bvalid;      // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_bvalid -> SMP_HPS:h2f_lw_BVALID
	wire   [2:0] smp_hps_h2f_lw_axi_master_awsize;      // SMP_HPS:h2f_lw_AWSIZE -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awsize
	wire         smp_hps_h2f_lw_axi_master_awvalid;     // SMP_HPS:h2f_lw_AWVALID -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_awvalid
	wire         smp_hps_h2f_lw_axi_master_rvalid;      // mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_rvalid -> SMP_HPS:h2f_lw_RVALID
	wire         mm_interconnect_0_pio_0_s1_chipselect; // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;   // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;    // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;      // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;  // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         rst_controller_reset_out_reset;        // rst_controller:reset_out -> [mm_interconnect_0:pio_0_reset_reset_bridge_in_reset_reset, pio_0:reset_n]
	wire         rst_controller_001_reset_out_reset;    // rst_controller_001:reset_out -> mm_interconnect_0:SMP_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	hps_design_SMP_HPS #(
		.F2S_Width (0),
		.S2F_Width (0)
	) smp_hps (
		.mem_a          (hps_ddr_mem_a),                     //            memory.mem_a
		.mem_ba         (hps_ddr_mem_ba),                    //                  .mem_ba
		.mem_ck         (hps_ddr_mem_ck),                    //                  .mem_ck
		.mem_ck_n       (hps_ddr_mem_ck_n),                  //                  .mem_ck_n
		.mem_cke        (hps_ddr_mem_cke),                   //                  .mem_cke
		.mem_cs_n       (hps_ddr_mem_cs_n),                  //                  .mem_cs_n
		.mem_ras_n      (hps_ddr_mem_ras_n),                 //                  .mem_ras_n
		.mem_cas_n      (hps_ddr_mem_cas_n),                 //                  .mem_cas_n
		.mem_we_n       (hps_ddr_mem_we_n),                  //                  .mem_we_n
		.mem_reset_n    (hps_ddr_mem_reset_n),               //                  .mem_reset_n
		.mem_dq         (hps_ddr_mem_dq),                    //                  .mem_dq
		.mem_dqs        (hps_ddr_mem_dqs),                   //                  .mem_dqs
		.mem_dqs_n      (hps_ddr_mem_dqs_n),                 //                  .mem_dqs_n
		.mem_odt        (hps_ddr_mem_odt),                   //                  .mem_odt
		.mem_dm         (hps_ddr_mem_dm),                    //                  .mem_dm
		.oct_rzqin      (hps_ddr_oct_rzqin),                 //                  .oct_rzqin
		.h2f_rst_n      (smp_hps_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_lw_axi_clk (pll_0_outclk0_clk),                 //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID    (smp_hps_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR  (smp_hps_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN   (smp_hps_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE  (smp_hps_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST (smp_hps_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK  (smp_hps_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE (smp_hps_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT  (smp_hps_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID (smp_hps_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY (smp_hps_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID     (smp_hps_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA   (smp_hps_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB   (smp_hps_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST   (smp_hps_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID  (smp_hps_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY  (smp_hps_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID     (smp_hps_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP   (smp_hps_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID  (smp_hps_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY  (smp_hps_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID    (smp_hps_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR  (smp_hps_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN   (smp_hps_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE  (smp_hps_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST (smp_hps_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK  (smp_hps_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE (smp_hps_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT  (smp_hps_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID (smp_hps_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY (smp_hps_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID     (smp_hps_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA   (smp_hps_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP   (smp_hps_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST   (smp_hps_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID  (smp_hps_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY  (smp_hps_h2f_lw_axi_master_rready)   //                  .rready
	);

	hps_design_pio_0 pio_0 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                            // external_connection.export
	);

	hps_design_pll_0 pll_0 (
		.refclk   (clk_clk),                  //  refclk.clk
		.rst      (~smp_hps_h2f_reset_reset), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),        // outclk0.clk
		.outclk_1 (),                         // outclk1.clk
		.outclk_2 (pll_0_sdram_clk),          // outclk2.clk
		.locked   ()                          // (terminated)
	);

	hps_design_mm_interconnect_0 mm_interconnect_0 (
		.SMP_HPS_h2f_lw_axi_master_awid                                        (smp_hps_h2f_lw_axi_master_awid),        //                                       SMP_HPS_h2f_lw_axi_master.awid
		.SMP_HPS_h2f_lw_axi_master_awaddr                                      (smp_hps_h2f_lw_axi_master_awaddr),      //                                                                .awaddr
		.SMP_HPS_h2f_lw_axi_master_awlen                                       (smp_hps_h2f_lw_axi_master_awlen),       //                                                                .awlen
		.SMP_HPS_h2f_lw_axi_master_awsize                                      (smp_hps_h2f_lw_axi_master_awsize),      //                                                                .awsize
		.SMP_HPS_h2f_lw_axi_master_awburst                                     (smp_hps_h2f_lw_axi_master_awburst),     //                                                                .awburst
		.SMP_HPS_h2f_lw_axi_master_awlock                                      (smp_hps_h2f_lw_axi_master_awlock),      //                                                                .awlock
		.SMP_HPS_h2f_lw_axi_master_awcache                                     (smp_hps_h2f_lw_axi_master_awcache),     //                                                                .awcache
		.SMP_HPS_h2f_lw_axi_master_awprot                                      (smp_hps_h2f_lw_axi_master_awprot),      //                                                                .awprot
		.SMP_HPS_h2f_lw_axi_master_awvalid                                     (smp_hps_h2f_lw_axi_master_awvalid),     //                                                                .awvalid
		.SMP_HPS_h2f_lw_axi_master_awready                                     (smp_hps_h2f_lw_axi_master_awready),     //                                                                .awready
		.SMP_HPS_h2f_lw_axi_master_wid                                         (smp_hps_h2f_lw_axi_master_wid),         //                                                                .wid
		.SMP_HPS_h2f_lw_axi_master_wdata                                       (smp_hps_h2f_lw_axi_master_wdata),       //                                                                .wdata
		.SMP_HPS_h2f_lw_axi_master_wstrb                                       (smp_hps_h2f_lw_axi_master_wstrb),       //                                                                .wstrb
		.SMP_HPS_h2f_lw_axi_master_wlast                                       (smp_hps_h2f_lw_axi_master_wlast),       //                                                                .wlast
		.SMP_HPS_h2f_lw_axi_master_wvalid                                      (smp_hps_h2f_lw_axi_master_wvalid),      //                                                                .wvalid
		.SMP_HPS_h2f_lw_axi_master_wready                                      (smp_hps_h2f_lw_axi_master_wready),      //                                                                .wready
		.SMP_HPS_h2f_lw_axi_master_bid                                         (smp_hps_h2f_lw_axi_master_bid),         //                                                                .bid
		.SMP_HPS_h2f_lw_axi_master_bresp                                       (smp_hps_h2f_lw_axi_master_bresp),       //                                                                .bresp
		.SMP_HPS_h2f_lw_axi_master_bvalid                                      (smp_hps_h2f_lw_axi_master_bvalid),      //                                                                .bvalid
		.SMP_HPS_h2f_lw_axi_master_bready                                      (smp_hps_h2f_lw_axi_master_bready),      //                                                                .bready
		.SMP_HPS_h2f_lw_axi_master_arid                                        (smp_hps_h2f_lw_axi_master_arid),        //                                                                .arid
		.SMP_HPS_h2f_lw_axi_master_araddr                                      (smp_hps_h2f_lw_axi_master_araddr),      //                                                                .araddr
		.SMP_HPS_h2f_lw_axi_master_arlen                                       (smp_hps_h2f_lw_axi_master_arlen),       //                                                                .arlen
		.SMP_HPS_h2f_lw_axi_master_arsize                                      (smp_hps_h2f_lw_axi_master_arsize),      //                                                                .arsize
		.SMP_HPS_h2f_lw_axi_master_arburst                                     (smp_hps_h2f_lw_axi_master_arburst),     //                                                                .arburst
		.SMP_HPS_h2f_lw_axi_master_arlock                                      (smp_hps_h2f_lw_axi_master_arlock),      //                                                                .arlock
		.SMP_HPS_h2f_lw_axi_master_arcache                                     (smp_hps_h2f_lw_axi_master_arcache),     //                                                                .arcache
		.SMP_HPS_h2f_lw_axi_master_arprot                                      (smp_hps_h2f_lw_axi_master_arprot),      //                                                                .arprot
		.SMP_HPS_h2f_lw_axi_master_arvalid                                     (smp_hps_h2f_lw_axi_master_arvalid),     //                                                                .arvalid
		.SMP_HPS_h2f_lw_axi_master_arready                                     (smp_hps_h2f_lw_axi_master_arready),     //                                                                .arready
		.SMP_HPS_h2f_lw_axi_master_rid                                         (smp_hps_h2f_lw_axi_master_rid),         //                                                                .rid
		.SMP_HPS_h2f_lw_axi_master_rdata                                       (smp_hps_h2f_lw_axi_master_rdata),       //                                                                .rdata
		.SMP_HPS_h2f_lw_axi_master_rresp                                       (smp_hps_h2f_lw_axi_master_rresp),       //                                                                .rresp
		.SMP_HPS_h2f_lw_axi_master_rlast                                       (smp_hps_h2f_lw_axi_master_rlast),       //                                                                .rlast
		.SMP_HPS_h2f_lw_axi_master_rvalid                                      (smp_hps_h2f_lw_axi_master_rvalid),      //                                                                .rvalid
		.SMP_HPS_h2f_lw_axi_master_rready                                      (smp_hps_h2f_lw_axi_master_rready),      //                                                                .rready
		.pll_0_outclk0_clk                                                     (pll_0_outclk0_clk),                     //                                                   pll_0_outclk0.clk
		.pio_0_reset_reset_bridge_in_reset_reset                               (rst_controller_reset_out_reset),        //                               pio_0_reset_reset_bridge_in_reset.reset
		.SMP_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),    // SMP_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.pio_0_s1_address                                                      (mm_interconnect_0_pio_0_s1_address),    //                                                        pio_0_s1.address
		.pio_0_s1_write                                                        (mm_interconnect_0_pio_0_s1_write),      //                                                                .write
		.pio_0_s1_readdata                                                     (mm_interconnect_0_pio_0_s1_readdata),   //                                                                .readdata
		.pio_0_s1_writedata                                                    (mm_interconnect_0_pio_0_s1_writedata),  //                                                                .writedata
		.pio_0_s1_chipselect                                                   (mm_interconnect_0_pio_0_s1_chipselect)  //                                                                .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~smp_hps_h2f_reset_reset),       // reset_in0.reset
		.clk            (pll_0_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~smp_hps_h2f_reset_reset),           // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
