// soc_design.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module soc_design (
		output wire [12:0] dram_addr,    //     dram.addr
		output wire [1:0]  dram_ba,      //         .ba
		output wire        dram_cas_n,   //         .cas_n
		output wire        dram_cke,     //         .cke
		output wire        dram_cs_n,    //         .cs_n
		inout  wire [15:0] dram_dq,      //         .dq
		output wire [1:0]  dram_dqm,     //         .dqm
		output wire        dram_ras_n,   //         .ras_n
		output wire        dram_we_n,    //         .we_n
		output wire        dram_clk_clk, // dram_clk.clk
		input  wire        fpga_reset_n, //     fpga.reset_n
		input  wire        ref_clk,      //      ref.clk
		input  wire        uart_RXD,     //     uart.RXD
		output wire        uart_TXD      //         .TXD
	);

	wire         system_pll_outclk0_clk;                                    // system_pll:outclk_0 -> [JTAG:clk, SDRAM:clk, SRAM:clk, Sys_Timer:clk, SystemID:clock, UART_COM:clk, irq_mapper:clk, mm_interconnect_0:system_pll_outclk0_clk, niosII_core:clk, rst_controller:clk]
	wire  [31:0] niosii_core_data_master_readdata;                          // mm_interconnect_0:niosII_core_data_master_readdata -> niosII_core:d_readdata
	wire         niosii_core_data_master_waitrequest;                       // mm_interconnect_0:niosII_core_data_master_waitrequest -> niosII_core:d_waitrequest
	wire         niosii_core_data_master_debugaccess;                       // niosII_core:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:niosII_core_data_master_debugaccess
	wire  [26:0] niosii_core_data_master_address;                           // niosII_core:d_address -> mm_interconnect_0:niosII_core_data_master_address
	wire   [3:0] niosii_core_data_master_byteenable;                        // niosII_core:d_byteenable -> mm_interconnect_0:niosII_core_data_master_byteenable
	wire         niosii_core_data_master_read;                              // niosII_core:d_read -> mm_interconnect_0:niosII_core_data_master_read
	wire         niosii_core_data_master_readdatavalid;                     // mm_interconnect_0:niosII_core_data_master_readdatavalid -> niosII_core:d_readdatavalid
	wire         niosii_core_data_master_write;                             // niosII_core:d_write -> mm_interconnect_0:niosII_core_data_master_write
	wire  [31:0] niosii_core_data_master_writedata;                         // niosII_core:d_writedata -> mm_interconnect_0:niosII_core_data_master_writedata
	wire   [3:0] niosii_core_data_master_burstcount;                        // niosII_core:d_burstcount -> mm_interconnect_0:niosII_core_data_master_burstcount
	wire  [31:0] niosii_core_instruction_master_readdata;                   // mm_interconnect_0:niosII_core_instruction_master_readdata -> niosII_core:i_readdata
	wire         niosii_core_instruction_master_waitrequest;                // mm_interconnect_0:niosII_core_instruction_master_waitrequest -> niosII_core:i_waitrequest
	wire  [26:0] niosii_core_instruction_master_address;                    // niosII_core:i_address -> mm_interconnect_0:niosII_core_instruction_master_address
	wire         niosii_core_instruction_master_read;                       // niosII_core:i_read -> mm_interconnect_0:niosII_core_instruction_master_read
	wire         niosii_core_instruction_master_readdatavalid;              // mm_interconnect_0:niosII_core_instruction_master_readdatavalid -> niosII_core:i_readdatavalid
	wire   [3:0] niosii_core_instruction_master_burstcount;                 // niosII_core:i_burstcount -> mm_interconnect_0:niosII_core_instruction_master_burstcount
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;       // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;         // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;      // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;          // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;             // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;            // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;        // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire         mm_interconnect_0_uart_com_avalon_rs232_slave_chipselect;  // mm_interconnect_0:UART_COM_avalon_rs232_slave_chipselect -> UART_COM:chipselect
	wire  [31:0] mm_interconnect_0_uart_com_avalon_rs232_slave_readdata;    // UART_COM:readdata -> mm_interconnect_0:UART_COM_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_uart_com_avalon_rs232_slave_address;     // mm_interconnect_0:UART_COM_avalon_rs232_slave_address -> UART_COM:address
	wire         mm_interconnect_0_uart_com_avalon_rs232_slave_read;        // mm_interconnect_0:UART_COM_avalon_rs232_slave_read -> UART_COM:read
	wire   [3:0] mm_interconnect_0_uart_com_avalon_rs232_slave_byteenable;  // mm_interconnect_0:UART_COM_avalon_rs232_slave_byteenable -> UART_COM:byteenable
	wire         mm_interconnect_0_uart_com_avalon_rs232_slave_write;       // mm_interconnect_0:UART_COM_avalon_rs232_slave_write -> UART_COM:write
	wire  [31:0] mm_interconnect_0_uart_com_avalon_rs232_slave_writedata;   // mm_interconnect_0:UART_COM_avalon_rs232_slave_writedata -> UART_COM:writedata
	wire  [31:0] mm_interconnect_0_systemid_control_slave_readdata;         // SystemID:readdata -> mm_interconnect_0:SystemID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_systemid_control_slave_address;          // mm_interconnect_0:SystemID_control_slave_address -> SystemID:address
	wire  [31:0] mm_interconnect_0_niosii_core_debug_mem_slave_readdata;    // niosII_core:debug_mem_slave_readdata -> mm_interconnect_0:niosII_core_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosii_core_debug_mem_slave_waitrequest; // niosII_core:debug_mem_slave_waitrequest -> mm_interconnect_0:niosII_core_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosii_core_debug_mem_slave_debugaccess; // mm_interconnect_0:niosII_core_debug_mem_slave_debugaccess -> niosII_core:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosii_core_debug_mem_slave_address;     // mm_interconnect_0:niosII_core_debug_mem_slave_address -> niosII_core:debug_mem_slave_address
	wire         mm_interconnect_0_niosii_core_debug_mem_slave_read;        // mm_interconnect_0:niosII_core_debug_mem_slave_read -> niosII_core:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosii_core_debug_mem_slave_byteenable;  // mm_interconnect_0:niosII_core_debug_mem_slave_byteenable -> niosII_core:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosii_core_debug_mem_slave_write;       // mm_interconnect_0:niosII_core_debug_mem_slave_write -> niosII_core:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosii_core_debug_mem_slave_writedata;   // mm_interconnect_0:niosII_core_debug_mem_slave_writedata -> niosII_core:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                      // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                        // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire  [14:0] mm_interconnect_0_sram_s1_address;                         // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                      // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                           // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                       // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                           // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         mm_interconnect_0_sys_timer_s1_chipselect;                 // mm_interconnect_0:Sys_Timer_s1_chipselect -> Sys_Timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_timer_s1_readdata;                   // Sys_Timer:readdata -> mm_interconnect_0:Sys_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_timer_s1_address;                    // mm_interconnect_0:Sys_Timer_s1_address -> Sys_Timer:address
	wire         mm_interconnect_0_sys_timer_s1_write;                      // mm_interconnect_0:Sys_Timer_s1_write -> Sys_Timer:write_n
	wire  [15:0] mm_interconnect_0_sys_timer_s1_writedata;                  // mm_interconnect_0:Sys_Timer_s1_writedata -> Sys_Timer:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         irq_mapper_receiver0_irq;                                  // UART_COM:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // JTAG:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // Sys_Timer:irq -> irq_mapper:receiver2_irq
	wire  [31:0] niosii_core_irq_irq;                                       // irq_mapper:sender_irq -> niosII_core:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [JTAG:rst_n, SDRAM:reset_n, SRAM:reset, Sys_Timer:reset_n, SystemID:reset_n, UART_COM:reset, irq_mapper:reset, mm_interconnect_0:niosII_core_reset_reset_bridge_in_reset_reset, niosII_core:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [SRAM:reset_req, niosII_core:reset_req, rst_translator:reset_req_in]

	soc_design_JTAG jtag (
		.clk            (system_pll_outclk0_clk),                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                              //               irq.irq
	);

	soc_design_SDRAM sdram (
		.clk            (system_pll_outclk0_clk),                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (dram_addr),                                //  wire.export
		.zs_ba          (dram_ba),                                  //      .export
		.zs_cas_n       (dram_cas_n),                               //      .export
		.zs_cke         (dram_cke),                                 //      .export
		.zs_cs_n        (dram_cs_n),                                //      .export
		.zs_dq          (dram_dq),                                  //      .export
		.zs_dqm         (dram_dqm),                                 //      .export
		.zs_ras_n       (dram_ras_n),                               //      .export
		.zs_we_n        (dram_we_n)                                 //      .export
	);

	soc_design_SRAM sram (
		.clk        (system_pll_outclk0_clk),               //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)    //       .reset_req
	);

	soc_design_Sys_Timer sys_timer (
		.clk        (system_pll_outclk0_clk),                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_sys_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                   //   irq.irq
	);

	soc_design_SystemID systemid (
		.clock    (system_pll_outclk0_clk),                            //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_systemid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_systemid_control_slave_address)   //              .address
	);

	soc_design_UART_COM uart_com (
		.clk        (system_pll_outclk0_clk),                                   //                clk.clk
		.reset      (rst_controller_reset_out_reset),                           //              reset.reset
		.address    (mm_interconnect_0_uart_com_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_uart_com_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_uart_com_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_uart_com_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_uart_com_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_uart_com_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_uart_com_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver0_irq),                                 //          interrupt.irq
		.UART_RXD   (uart_RXD),                                                 // external_interface.export
		.UART_TXD   (uart_TXD)                                                  //                   .export
	);

	soc_design_niosII_core niosii_core (
		.clk                                 (system_pll_outclk0_clk),                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                           //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                        //                          .reset_req
		.d_address                           (niosii_core_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosii_core_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosii_core_data_master_read),                              //                          .read
		.d_readdata                          (niosii_core_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosii_core_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosii_core_data_master_write),                             //                          .write
		.d_writedata                         (niosii_core_data_master_writedata),                         //                          .writedata
		.d_burstcount                        (niosii_core_data_master_burstcount),                        //                          .burstcount
		.d_readdatavalid                     (niosii_core_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (niosii_core_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosii_core_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosii_core_instruction_master_read),                       //                          .read
		.i_readdata                          (niosii_core_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosii_core_instruction_master_waitrequest),                //                          .waitrequest
		.i_burstcount                        (niosii_core_instruction_master_burstcount),                 //                          .burstcount
		.i_readdatavalid                     (niosii_core_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (niosii_core_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                          //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosii_core_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosii_core_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosii_core_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosii_core_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosii_core_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosii_core_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosii_core_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosii_core_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                           // custom_instruction_master.readra
	);

	soc_design_system_pll system_pll (
		.refclk   (ref_clk),                //  refclk.clk
		.rst      (~fpga_reset_n),          //   reset.reset
		.outclk_0 (system_pll_outclk0_clk), // outclk0.clk
		.outclk_1 (dram_clk_clk),           // outclk1.clk
		.locked   ()                        // (terminated)
	);

	soc_design_mm_interconnect_0 mm_interconnect_0 (
		.system_pll_outclk0_clk                        (system_pll_outclk0_clk),                                    //                      system_pll_outclk0.clk
		.niosII_core_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // niosII_core_reset_reset_bridge_in_reset.reset
		.niosII_core_data_master_address               (niosii_core_data_master_address),                           //                 niosII_core_data_master.address
		.niosII_core_data_master_waitrequest           (niosii_core_data_master_waitrequest),                       //                                        .waitrequest
		.niosII_core_data_master_burstcount            (niosii_core_data_master_burstcount),                        //                                        .burstcount
		.niosII_core_data_master_byteenable            (niosii_core_data_master_byteenable),                        //                                        .byteenable
		.niosII_core_data_master_read                  (niosii_core_data_master_read),                              //                                        .read
		.niosII_core_data_master_readdata              (niosii_core_data_master_readdata),                          //                                        .readdata
		.niosII_core_data_master_readdatavalid         (niosii_core_data_master_readdatavalid),                     //                                        .readdatavalid
		.niosII_core_data_master_write                 (niosii_core_data_master_write),                             //                                        .write
		.niosII_core_data_master_writedata             (niosii_core_data_master_writedata),                         //                                        .writedata
		.niosII_core_data_master_debugaccess           (niosii_core_data_master_debugaccess),                       //                                        .debugaccess
		.niosII_core_instruction_master_address        (niosii_core_instruction_master_address),                    //          niosII_core_instruction_master.address
		.niosII_core_instruction_master_waitrequest    (niosii_core_instruction_master_waitrequest),                //                                        .waitrequest
		.niosII_core_instruction_master_burstcount     (niosii_core_instruction_master_burstcount),                 //                                        .burstcount
		.niosII_core_instruction_master_read           (niosii_core_instruction_master_read),                       //                                        .read
		.niosII_core_instruction_master_readdata       (niosii_core_instruction_master_readdata),                   //                                        .readdata
		.niosII_core_instruction_master_readdatavalid  (niosii_core_instruction_master_readdatavalid),              //                                        .readdatavalid
		.JTAG_avalon_jtag_slave_address                (mm_interconnect_0_jtag_avalon_jtag_slave_address),          //                  JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_avalon_jtag_slave_write),            //                                        .write
		.JTAG_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_avalon_jtag_slave_read),             //                                        .read
		.JTAG_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),         //                                        .readdata
		.JTAG_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),        //                                        .writedata
		.JTAG_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),      //                                        .waitrequest
		.JTAG_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),       //                                        .chipselect
		.niosII_core_debug_mem_slave_address           (mm_interconnect_0_niosii_core_debug_mem_slave_address),     //             niosII_core_debug_mem_slave.address
		.niosII_core_debug_mem_slave_write             (mm_interconnect_0_niosii_core_debug_mem_slave_write),       //                                        .write
		.niosII_core_debug_mem_slave_read              (mm_interconnect_0_niosii_core_debug_mem_slave_read),        //                                        .read
		.niosII_core_debug_mem_slave_readdata          (mm_interconnect_0_niosii_core_debug_mem_slave_readdata),    //                                        .readdata
		.niosII_core_debug_mem_slave_writedata         (mm_interconnect_0_niosii_core_debug_mem_slave_writedata),   //                                        .writedata
		.niosII_core_debug_mem_slave_byteenable        (mm_interconnect_0_niosii_core_debug_mem_slave_byteenable),  //                                        .byteenable
		.niosII_core_debug_mem_slave_waitrequest       (mm_interconnect_0_niosii_core_debug_mem_slave_waitrequest), //                                        .waitrequest
		.niosII_core_debug_mem_slave_debugaccess       (mm_interconnect_0_niosii_core_debug_mem_slave_debugaccess), //                                        .debugaccess
		.SDRAM_s1_address                              (mm_interconnect_0_sdram_s1_address),                        //                                SDRAM_s1.address
		.SDRAM_s1_write                                (mm_interconnect_0_sdram_s1_write),                          //                                        .write
		.SDRAM_s1_read                                 (mm_interconnect_0_sdram_s1_read),                           //                                        .read
		.SDRAM_s1_readdata                             (mm_interconnect_0_sdram_s1_readdata),                       //                                        .readdata
		.SDRAM_s1_writedata                            (mm_interconnect_0_sdram_s1_writedata),                      //                                        .writedata
		.SDRAM_s1_byteenable                           (mm_interconnect_0_sdram_s1_byteenable),                     //                                        .byteenable
		.SDRAM_s1_readdatavalid                        (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                        .readdatavalid
		.SDRAM_s1_waitrequest                          (mm_interconnect_0_sdram_s1_waitrequest),                    //                                        .waitrequest
		.SDRAM_s1_chipselect                           (mm_interconnect_0_sdram_s1_chipselect),                     //                                        .chipselect
		.SRAM_s1_address                               (mm_interconnect_0_sram_s1_address),                         //                                 SRAM_s1.address
		.SRAM_s1_write                                 (mm_interconnect_0_sram_s1_write),                           //                                        .write
		.SRAM_s1_readdata                              (mm_interconnect_0_sram_s1_readdata),                        //                                        .readdata
		.SRAM_s1_writedata                             (mm_interconnect_0_sram_s1_writedata),                       //                                        .writedata
		.SRAM_s1_byteenable                            (mm_interconnect_0_sram_s1_byteenable),                      //                                        .byteenable
		.SRAM_s1_chipselect                            (mm_interconnect_0_sram_s1_chipselect),                      //                                        .chipselect
		.SRAM_s1_clken                                 (mm_interconnect_0_sram_s1_clken),                           //                                        .clken
		.Sys_Timer_s1_address                          (mm_interconnect_0_sys_timer_s1_address),                    //                            Sys_Timer_s1.address
		.Sys_Timer_s1_write                            (mm_interconnect_0_sys_timer_s1_write),                      //                                        .write
		.Sys_Timer_s1_readdata                         (mm_interconnect_0_sys_timer_s1_readdata),                   //                                        .readdata
		.Sys_Timer_s1_writedata                        (mm_interconnect_0_sys_timer_s1_writedata),                  //                                        .writedata
		.Sys_Timer_s1_chipselect                       (mm_interconnect_0_sys_timer_s1_chipselect),                 //                                        .chipselect
		.SystemID_control_slave_address                (mm_interconnect_0_systemid_control_slave_address),          //                  SystemID_control_slave.address
		.SystemID_control_slave_readdata               (mm_interconnect_0_systemid_control_slave_readdata),         //                                        .readdata
		.UART_COM_avalon_rs232_slave_address           (mm_interconnect_0_uart_com_avalon_rs232_slave_address),     //             UART_COM_avalon_rs232_slave.address
		.UART_COM_avalon_rs232_slave_write             (mm_interconnect_0_uart_com_avalon_rs232_slave_write),       //                                        .write
		.UART_COM_avalon_rs232_slave_read              (mm_interconnect_0_uart_com_avalon_rs232_slave_read),        //                                        .read
		.UART_COM_avalon_rs232_slave_readdata          (mm_interconnect_0_uart_com_avalon_rs232_slave_readdata),    //                                        .readdata
		.UART_COM_avalon_rs232_slave_writedata         (mm_interconnect_0_uart_com_avalon_rs232_slave_writedata),   //                                        .writedata
		.UART_COM_avalon_rs232_slave_byteenable        (mm_interconnect_0_uart_com_avalon_rs232_slave_byteenable),  //                                        .byteenable
		.UART_COM_avalon_rs232_slave_chipselect        (mm_interconnect_0_uart_com_avalon_rs232_slave_chipselect)   //                                        .chipselect
	);

	soc_design_irq_mapper irq_mapper (
		.clk           (system_pll_outclk0_clk),         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (niosii_core_irq_irq)             //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~fpga_reset_n),                      // reset_in0.reset
		.clk            (system_pll_outclk0_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
